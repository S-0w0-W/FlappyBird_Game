LIBRARY IEEE;
USE  IEEE.STD_LOGIC_1164.all;
USE  IEEE.STD_LOGIC_UNSIGNED.all;
use ieee.numeric_std.all;

ENTITY pipeDrawer IS
	GENERIC(
		PIPE_WIDTH 					: INTEGER RANGE 0 TO 100 := 60;
		PIPE_GAP 					: INTEGER RANGE 0 TO 300 := 150;
		PIPE_LIP_HEIGHT			: INTEGER RANGE 0 TO 100 := 40;
		PIPE_LIP_EDGE				: INTEGER RANGE 0 TO 10 := 4;
		
		highLightIn 				: integer range 0 to 40 := 16;
		highLightOut 				: integer range 0 to 40 := 27;
		midToneIn					: integer range 0 to 40 := 8;
		midToneOut 					: integer range 0 to 40 := 40
		
	);
	
	PORT(
		clk25MHz, vertSync		: IN	STD_LOGIC;
		pipeY, pipeX				: IN	SIGNED(10 DOWNTO 0);
		pixel_row, pixel_col		: IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		
		R, G, B						: OUT	STD_LOGIC_VECTOR(3 DOWNTO 0);
		A								: OUT	STD_LOGIC
		
	);
END ENTITY pipeDrawer;

architecture drawBehaviour OF pipeDrawer IS
	SIGNAL pipeOn : STD_LOGIC;
	SIGNAL colour : STD_LOGIC_VECTOR(1 DOWNTO 0);
	SIGNAL prevPipeX, prevPipeY : SIGNED(10 DOWNTO 0);
begin
	--	
	A <= pipeOn;
	R <= "0010" when colour = "00" ELSE
		  "0010" when colour = "01" ELSE
		  "0010" when colour = "10" ELSE
		  "0000";
		  
	G <= "1111" when colour = "00" ELSE
		  "1010" when colour = "01" ELSE
		  "0111" when colour = "10" ELSE
		  "0000";
		  
	B <= "0010" when colour = "00" ELSE
		  "0010" when colour = "01" ELSE
		  "0010" when colour = "10" ELSE
		  "0000";
	--pipe
	pipeGen : PROCESS(pixel_row, pixel_col, prevPipeX, prevPipeY)
	BEGin
		IF (signed('0' & pixel_row) <= prevPipeY - to_signed(2, prevPipeY'length)) and 
			(signed('0' & pixel_row) >= prevPipeY - to_signed(PIPE_GAP - 2, prevPipeY'length)) THEN
			pipeOn <= '0';
		
		ELSIF (signed('0' & pixel_row) <= prevPipeY) and 
				(signed('0' & pixel_row) >= prevPipeY - to_signed(PIPE_GAP, prevPipeY'length)) and
				(signed('0' & pixel_col) <= prevPipeX) and 
				(signed('0' & pixel_col) >= prevPipeX - to_signed(PIPE_WIDTH, prevPipeY'length))	THEN
				pipeOn <= '1';
				colour <= "11";
				
		ELSIF (signed('0' & pixel_row) <= prevPipeY + to_signed(PIPE_LIP_HEIGHT - 2, prevPipeY'length)) and 
				(signed('0' & pixel_row) >= prevPipeY - to_signed(PIPE_GAP + PIPE_LIP_HEIGHT - 2, prevPipeY'length)) THEN
			
			pipeOn <= '1';
			--HighLights of the smaller pipe
			IF (signed('0' & pixel_col) <= prevPipeX - to_signed(highLightIn, prevPipeX'length)) and 
				(signed('0' & pixel_col) >= prevPipeX - to_signed(highLightOut, prevPipeX'length)) THEN 
				colour <= "00"; 
				
			ELSIF (signed('0' & pixel_col) <= prevPipeX - to_signed(midToneIn, prevPipeX'length)) and 
					(signed('0' & pixel_col) >= prevPipeX - to_signed(midToneOut, prevPipeX'length)) THEN 
				colour <= "01"; 
			
			ELSIF (signed('0' & pixel_col) <= prevPipeX - to_signed(2, prevPipeY'length)) and 
					(signed('0' & pixel_col) >= prevPipeX - to_signed(PIPE_WIDTH - 2, prevPipeX'length)) THEN 
				colour <= "10";
			ELSIF (signed('0' & pixel_col) <= prevPipeX) and 
					(signed('0' & pixel_col) >= prevPipeX - to_signed(PIPE_WIDTH, prevPipeY'length)) THEN 
				colour <= "11"; 	
			ELSE
				pipeOn <= '0'; 
			END IF;
		ELSIF (signed('0' & pixel_row) <= prevPipeY + to_signed(PIPE_LIP_HEIGHT, prevPipeY'length)) and 
				(signed('0' & pixel_row) >= prevPipeY - to_signed(PIPE_GAP + PIPE_LIP_HEIGHT, prevPipeY'length)) and
				(signed('0' & pixel_col) <= prevPipeX) and 
				(signed('0' & pixel_col) >= prevPipeX - to_signed(PIPE_WIDTH, prevPipeY'length))	THEN
				pipeOn <= '1';
				colour <= "11";
		ELSE
			pipeOn <= '1';
			
			--HighLights of the smaller pipe
			IF (signed('0' & pixel_col) <= prevPipeX - to_signed(highLightIn + PIPE_LIP_EDGE, prevPipeY'length)) and 
				(signed('0' & pixel_col) >= prevPipeX - to_signed(highLightOut + PIPE_LIP_EDGE, prevPipeY'length)) THEN 
				colour <= "00"; 
				
			ELSIF (signed('0' & pixel_col) <= prevPipeX - to_signed(midToneIn + PIPE_LIP_EDGE, prevPipeY'length)) and 
					(signed('0' & pixel_col) >= prevPipeX - to_signed(midToneOut + PIPE_LIP_EDGE, prevPipeY'length)) THEN 
				colour <= "01"; 
			
			ELSIF (signed('0' & pixel_col) <= prevPipeX - to_signed(PIPE_LIP_EDGE + 2, prevPipeY'length)) and 
					(signed('0' & pixel_col) >= prevPipeX - to_signed(PIPE_WIDTH - PIPE_LIP_EDGE - 2, prevPipeY'length)) THEN 
				colour <= "10"; 
			
			ELSIF (signed('0' & pixel_col) <= prevPipeX - to_signed(PIPE_LIP_EDGE, prevPipeY'length)) and 
					(signed('0' & pixel_col) >= prevPipeX - to_signed(PIPE_WIDTH-PIPE_LIP_EDGE, prevPipeY'length)) THEN 
				colour <= "11"; 
			
			ELSE
				pipeOn <= '0'; 
			END IF; 
		END IF; 
	END PROCESS pipeGen; 
	
	--vertSync
	vert : PROCESS(clk25MHz)
	variable prevVert : STD_LOGIC := '0';
	BEGIn
		IF rising_edge(clk25MHz) THEN
			IF prevVert /= vertSync THEN
				prevVert := vertSync;
				prevPipeX <= pipeX;
				prevPipeY <= pipeY;
			ELSE
				prevVert := vertSync;
			END IF;
		END IF;
	
	END PROCESS vert;
end architecture drawBehaviour;